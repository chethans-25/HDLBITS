module top_module ( input a, input b, output out );
//mod_a is already available
  mod_a mod_a_i1 (.in1(a),.in2(b),.out(out));
endmodule
