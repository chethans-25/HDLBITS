module top_module(
  input clk,
  input in,
  input reset,
  output out);

	parameter A = 0, B = 1, C = 2, D = 3;
	reg [1:0] state, next_state;

  // State transition logic
	always @( * )
	begin
		case (state)
			A: next_state = in? B : A;
			B,D: next_state = in? B : C;
			C: next_state = in? D : A;
			default: next_state = state;
		endcase
	end
  
	// State flip-flops with asynchronous reset
	always @(posedge clk)
	begin
		state <= reset ? A : next_state;
	end
  
	// Output logic
	assign out = (state == D);

endmodule
